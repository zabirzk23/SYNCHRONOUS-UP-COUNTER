library verilog;
use verilog.vl_types.all;
entity UPCOUNTER_vlg_vec_tst is
end UPCOUNTER_vlg_vec_tst;
